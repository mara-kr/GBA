
module priority_eval (
    [19:0] BG,
    [19:0] OBJ);


endmodule priority_eval

/**lib - not sure if we want a separate file for this*/



