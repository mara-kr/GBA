/*module mixer ( input logic system_clock,
               input logic reset,
               input logic [23:0] channel1,
               input logic [23:0] channel2,
               input logic [23:0] channel3,
               input logic [23:0] channel4,
               input logic NR50,
               input logic NR51,
               output logic [23:0] output_wave_left,
               output logic [23:0] output_wave_right);

                //channel >> (master_volume << 1)
                
               always_comb begin
                         
               end
    
endmodule: mixer

*/