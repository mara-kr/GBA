`default_nettype none

module obj_register #(parameter WIDTH = 8) (
    input  logic clock, reset,
    output logic [WIDTH-1:0] q,
    input  logic [WIDTH-1:0] d,
    input  logic en, clear);

    always_ff @(posedge clock, negedge reset) begin
        if (reset) q <= {WIDTH{1'b0}};
        else if (clear) q <= {WIDTH{1'b0}};
        else if (en) q <= d;
    end
endmodule: obj_register

module obj_counter #(parameter WIDTH = 8) (
    input  logic clock, reset,
    output logic [WIDTH-1:0] q,
    input  logic en, clear);

    always_ff @(posedge clock, negedge reset) begin
        if (reset) q <= {WIDTH{1'b0}};
        else if (clear) q <= {WIDTH{1'b0}};
        else if (en) q <= q + 1;
    end
endmodule: obj_counter

module is_transparent (
    output logic        transparent,
    input  logic [15:0] data,
    input  logic        palettemode);

    assign transparent = (palettemode) ? |data[7:0] : |data[3:0];
endmodule: is_transparent

module within_preimage_checker (
    output logic        valid,
    input  logic [10:0] X, Y, hsize, vsize);

    assign valid = (X < hsize) & (Y < vsize);

endmodule: within_preimage_checker

module obj_data_unit (
    output logic  [7:0] palette_info,
    input  logic [15:0] data,
    input  logic [10:0] X,
    input  logic  [7:0] addr,
    input  logic  [3:0] palette_no,
    input  logic        palettemode);

    logic [7:0] data8;
    assign data8 = (addr[0]) ? data[15:8] : data[7:0];

    assign palette_info = (palettemode) ? data8 :
                    (X[0] ? {palette_no, data8[7:4]} : {palette_no, data[3:0]});

endmodule: obj_data_unit

module row_visible_unit (
    output logic       visible,
    input  logic [7:0] row, objy,
    input  logic [6:0] vsize,
    input  logic       rotation);

    logic [7:0] lowerbound;
    logic [7:0] adjust_objy;

    assign lowerbound = rotation ? objy - {2'b0, vsize} : objy;
    assign upperbound = lowerbound + {1'b0, vsize};
    assign visible = (row < upperbound) & (lowerbound[7] | (lowerbound <= row));

endmodule: row_visible_unit
